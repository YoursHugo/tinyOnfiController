module set_feature();
  onfi_cen=0;
end module